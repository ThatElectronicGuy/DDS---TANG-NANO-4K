Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.counter_8bit;
use work.counter_32bit;
use work.LSB_8bit_Shift_Register;
use work.LSB_32bit_Shift_Register;

entity top is
    Port (
            CLK_27MHZ : in STD_LOGIC;
            CLK_594MHZ : out STD_LOGIC;
            LED : out STD_LOGIC;
            CS32 : in STD_LOGIC;
            CS8 : in STD_LOGIC;
            MOSI : in STD_LOGIC;
            MSCLK : in STD_LOGIC -- MSCLK from uC side
         );
end top;

architecture Behavioral of top is

    -- internal signal clock generated by PLL
    signal clock_594MHZ : STD_LOGIC;
    --
    --
    constant MAX32 : unsigned (31 downto 0) := (others => '1');
    signal Q2 : STD_LOGIC_VECTOR (31 downto 0) := (others => '0');
    signal Q : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
    signal slow_clk : STD_LOGIC := '0';
    signal clk_div : unsigned (23 downto 0) := (others => '0');
    signal enableV : STD_LOGiC := '1';
    signal resetV : STD_LOGIC := '0';
    signal aresetV : STD_LOGIC := '0';
    signal LED_flag : STD_LOGIC := '0';
    --


    -- Signals necessary for Input demultiplexer
    signal Output32SPIIN : STD_LOGIC := '0';
    signal Output8SPIIN : STD_LOGIC := '0';
    signal Input_SPI : STD_LOGIC := '0';
    --

    -- Signals responsible for bit shift registers
    signal Q8BS : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
    signal Q32BS : STD_LOGIC_VECTOR (32 downto 0) := (others => '0');
    signal Reset_All : STD_LOGIC := '0';
    --------------------------------------------
begin

    -- Demultiplexer for SPI input
    Output32SPIIN <= Input_SPI when (CS32 = '0' and CS8 = '1') else '0';
    Output8SPIIN <= Input_SPI when (CS8 = '0' and CS32 = '1') else '0';
    --

    -- instantiating 8 bit shift register
    bit_shift_register_8 : entity work.LSB_8bit_Shift_Register
    port map
    (
        D => Output8,
        Q => Q8BS,
        CLK => MSCLK,
        RESET => Reset_All,
        ENABLE => not CS8
    );
    --

    -- instatiating 32 bit shift register
    bit_shift_register_32 : entity work.LSB_32bit_Shift_Register
    port map
    (
        D => Output32,
        Q => Q32BS,
        CLK => MSCLK,
        RESET => Reset_All,
        Enable => not CS32
    );
    --

    -- 





















-----------------------------------------------------------------------------------------------
    --instantiating 594 mhz clock pll entity
    PLL : entity work.Gowin_PLLVR
    port map
    (
        clkin => CLK_27MHZ,
        clkout => clock_594MHZ
    );


    --giving internal pll clock on output pin
    CLK_594MHZ <= clock_594MHZ;


    --
    process(CLK_27MHZ)      --      process of clock divider
    begin
        if rising_edge(CLK_27MHZ) then
        clk_div <= clk_div + 1;
        if clk_div = 135000 then
        slow_clk <= not slow_clk;
        clk_div <= (others => '0');
        end if;
        end if;
    end process;


    --
    --instantiating 8 bit counter
    LED_counter : entity work.counter_8bit
    port map (
        CLK => slow_clk,
        ENABLE => enableV,
        RESET => resetV,
        ARESET => aresetV,
        D => "00000001",
        Q => Q
    );
     


end Behavioral;