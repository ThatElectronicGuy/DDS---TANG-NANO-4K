Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.counter_8bit;
use work.counter_32bit;

entity top is
    Port (
            CLK_27MHZ : in STD_LOGIC;
            CLK_594MHZ : out STD_LOGIC;
            enable : in STD_LOGIC;
            RESET : in STD_LOGIC;
            ARESET : in STD_LOGIC;
            LED : out STD_LOGIC;
            debug_out : out STD_LOGIC;
            debug_PLL_594MHZ : out STD_LOGIC
         );
end top;

architecture Behavioral of top is

    -- internal signal clock generated by PLL
    signal clock_594MHZ : STD_LOGIC;
    --
    attribute syn_keep : boolean;    

    -- test signals
    signal Q2 : STD_LOGIC_VECTOR (31 downto 0) := (others => '0');
    signal Q : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
    constant MAX32 : unsigned (31 downto 0) := (others => '1');
    signal debug_PLL_594MHZ_s : STD_LOGIC := '0';
    attribute syn_keep of debug_PLL_594MHZ_s : signal is true;


    -- creating internal signal for oscillscope purposes
    signal internal_clock_27Mhz : STD_LOGIC;
    signal test_bit : STD_LOGIC := '0';
    attribute syn_keep of test_bit : signal is true;
    --

    --
    signal slow_clk : STD_LOGIC := '0';
    signal clk_div : unsigned (23 downto 0) := (others => '0');
    signal LED_flag : STD_LOGIC := '0';
    attribute syn_keep of LED_flag : signal is true;
    signal enableV : STD_LOGiC := '1';
    signal resetV : STD_LOGIC := '0';
    signal aresetV : STD_LOGIC := '0';
    --

begin
    
    --instantiating 594 mhz clock pll entity
    PLL : entity work.Gowin_PLLVR
    port map
    (
        clkin => CLK_27MHZ,
        clkout => clock_594MHZ
    );
    --giving internal pll clock on output pin
    CLK_594MHZ <= clock_594MHZ;

    --PLL 594 MHZ clock test
    PLL_clock_test : entity work.counter_32bit
    port map
    (
        CLK => clock_594MHZ,
        ENABLE => enableV,
        RESET => resetV,
        ARESET => aresetV,
        D => x"FFFFFFF1",
        Q => Q2
    );
    process (clock_594MHZ)
    begin
        enableV <= '1';
        if rising_edge(clock_594MHZ) then
        if unsigned(Q2) =  MAX32 then
        debug_PLL_594MHZ_s <= not debug_PLL_594MHZ_s;
        end if;
        end if;
        
    end process;

    debug_PLL_594MHZ <= debug_PLL_594MHZ_s;

    --
    




    internal_clock_27Mhz <= CLK_27MHZ;

    --create any process just to not have this signal ruled out by hidden processes
    process(internal_clock_27Mhz)
    begin
        if rising_edge(internal_clock_27Mhz) then
        test_bit <= not test_bit;
        end if;
    end process;
    debug_out <= test_bit;



    --
    process(CLK_27MHZ)      --      process of clock divider
    begin
        if rising_edge(CLK_27MHZ) then
        clk_div <= clk_div + 1;
        if clk_div = 135000 then
        slow_clk <= not slow_clk;
        clk_div <= (others => '0');
        end if;
        end if;
    end process;


    --
    --instantiating 8 bit counter
    LED_counter : entity work.counter_8bit
    port map (
        CLK => slow_clk,
        ENABLE => enableV,
        RESET => resetV,
        ARESET => aresetV,
        D => "00000001",
        Q => Q
    );
     
    process(slow_clk)
    begin
        enableV <= '1';
        if rising_edge(slow_clk) then
        if Q = "01111111" then
        LED_flag <= not LED_flag;
        resetV <= '1';
        else
        resetV <= '0';
        end if;
        end if;
    end process;

    LED <= LED_flag;

end Behavioral;